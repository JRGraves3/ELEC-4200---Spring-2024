`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/25/2024 11:27:57 AM
// Design Name: 
// Module Name: lab2_task4_part2
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lab2_task4_part2(
    input [3:0] a, b,
    input cin,
    output [3:0] s,
    output cout
    );
    
    wire w1, w2, w3;
    
    
endmodule
